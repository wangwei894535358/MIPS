`timescale 1ns / 1ps
module InstructionMem(instruction,address);
input[31:0] address;
output reg [31:0] instruction;
reg[31:0] Imemory[63:0];

integer k;

initial begin
	for(k=0;k<64;k=k+1)begin
		Imemory[k] = 32'b0;
	end
	//You can give your own code block here.
	//$t0: 01000 8, $t1: 01001: 9, $s0: 10000 16, $s1: 10001 17, $s2 10010 18 $s3 10011 19
	//
		 Imemory[0]  = 32'b10001100000100000000000000000000; 
		 Imemory[1]  = 32'b00000000000100000100000000100000; 
		 Imemory[2]  = 32'b00000000000100000100100000100000; 
		 Imemory[3]  = 32'b00000000000100000101000000100000;
		 Imemory[4]  = 32'b00010001000010010000000000000010;
		 Imemory[5]  = 32'b00000000000100001000100000100000;
		 Imemory[6]  = 32'b00000010001100001000100000100000;
		 Imemory[7]  = 32'b00000001000100000100000000100000;
		 Imemory[8]  = 32'b00000001010100000101000000100000;
		 Imemory[9]  = 32'b00000001001100000100100000100000;
		Imemory[10]  = 32'b00010001000010010000000000000010;
		Imemory[11]  = 32'b00000010001100001000100000100000;
		Imemory[12]  = 32'b00000010001100001000100000100000;
		Imemory[13]  = 32'b00000001001100000100100000100000;
		Imemory[14]  = 32'b10001100000010000000000000001000;
		Imemory[15]  = 32'b00000001010100000101000000100000;
		Imemory[16]  = 32'b00010001000010010000000000000010;
		Imemory[17]  = 32'b00000010001100001000100000100000;
		Imemory[18]  = 32'b00000010001100001000100000100000;
		Imemory[19]  = 32'b00000001001100000100100000100000;
		Imemory[20]  = 32'b00000001010100000101000000100000;
		Imemory[21]  = 32'b10001100000010000000000000001100;
		Imemory[22]  = 32'b00010001000010010000000000000010;
		Imemory[23]  = 32'b00000010001100001000100000100000;
		Imemory[24]  = 32'b00000010001100001000100000100000;
		Imemory[25]  = 32'b00000001000100000100000000100000;
		Imemory[26]  = 32'b00000001001100000100100000100000;
		Imemory[27]  = 32'b00010001000010010000000000000010;
		Imemory[28]  = 32'b00000010001100001000100000100000;
		Imemory[29]  = 32'b00000010001100001000100000100000;
		Imemory[30]  = 32'b10001100000010000000000000000000;
		Imemory[31]  = 32'b10001100000010010000000000000000;
		Imemory[32]  = 32'b00010001000010010000000000000010;
		Imemory[33]  = 32'b00000010001100001000100000100000;
		Imemory[34]  = 32'b00000010001100001000100000100000;
		Imemory[35]  = 32'b00000000000100000110000000100000;
		
		
		
		
		
		
		
	
	
		
	// lw $16, 0($0)  
	// add $8, $0, $16  
	// add $9, $0, $16  
	// add $10, $0, $16  
	// beq $8, $9, test2 
	// add $17, $0, $16	
	// add $17, $17, $16	
	// add $8, $8, $16	
	// add $10, $10, $16 	
	// add $9, $9, $16	
	// beq $8, $9, test3 
	// add $17, $17, $16	
	// add $17, $17, $16	
	// add $9, $9, $16	
	// lw $8, 8($0) 		
	// add $10, $10, $16 	
	// beq $8, $9, test4 
	// add $17, $17, $16 	
	// add $17, $17, $16	
	// add $9, $9, $16 	
	// add $10, $10, $16 	
	// lw $8, 12($0) 		
	// beq $8, $9, test5 
	// add $17, $17, $16 	
	// add $17, $17, $16 	
	// add $8, $8, $16 	
	// add $9, $9, $16   
	// beq $8, $9, test6 
	// add $17, $17, $16 	
	// add $17, $17, $16	
	// lw $8, 0($0) 		
	// lw $9, 0($0) 		
	// beq $8, $9, test7	
	// add $17, $17, $16	
	// add $17, $17, $16	
	// add $12, $0, $16 		

end

always @ (address)
	begin
		instruction <= Imemory[address[13:2]];
end
endmodule
